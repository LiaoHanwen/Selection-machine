--------------------------------------------------------------------------------
--save music
--
--input clock enable
--output tone
--
--integration test 10.31
--------------------------------------------------------------------------------

--------------------------------------------------------------------------------
--head

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

--head
--------------------------------------------------------------------------------


--------------------------------------------------------------------------------
--entity

entity save_music is
  port (
  	--in
	clock:in std_logic;
	enable:in std_logic;

	--out
	tone:out std_logic_vector(15 downto 0)
  ) ;
end entity ; -- save_music

--entity
--------------------------------------------------------------------------------

--------------------------------------------------------------------------------
--architecture

architecture arch of save_music is
	----------------------------------------------------------------------------
	--signal

	signal count: integer range 0 to 64 :=0;

	--signal
	----------------------------------------------------------------------------

begin

	----------------------------------------------------------------------------
	--play

	play : process( clock )
	begin
		if enable = '1' then
			if clock'event and clock='1' then
				if count < 61 then                             
					case count is                                 
						when 0 => tone <=b"0000000000000100";
						when 1 => tone <=b"0000000000001000";
						when 2 => tone <=b"0000000000010000";
						when 3 => tone <=b"0000000000001000";
						when 4 => tone <=b"0000000000000100";
						when 5 => tone <=b"0000000000001000";
						when 6 => tone <=b"0000000000010000";
						when 7 => tone <=b"0000000000001000";
						when 8 => tone <=b"0000000000000100";
						when 9 => tone <=b"0000000000001000";
						when 10 => tone <=b"0000000000010000";
						when 11 => tone <=b"0000000000010000";
						when 12 => tone <=b"0000000000001000";
						when 13 => tone <=b"0000000000010000";
						when 14 => tone <=b"0000010000000000";
						when 15 => tone <=b"0000000100000000";
						when 16 => tone <=b"0000000100000000";
						when 17 => tone <=b"0000000000000010";
						when 18 => tone <=b"0000000000000100";
						when 19 => tone <=b"0000000000001000";
						when 20 => tone <=b"0000000000000100";
						when 21 => tone <=b"0000000000001000";
						when 22 => tone <=b"0000001000000000";
						when 23 => tone <=b"0000000001000000";
						when 24 => tone <=b"0000000001000000";
						when 25 => tone <=b"0000000000000010";
						when 26 => tone <=b"0000000000000100";
						when 27 => tone <=b"0000000000001000";
						when 28 => tone <=b"0000000000000100";
						when 29 => tone <=b"0000000000001000";
						when 30 => tone <=b"0000000000100000";
						when 31 => tone <=b"0000000000010000";
						when 32 => tone <=b"0000000000010000";
						when 33 => tone <=b"0000000000000100";
						when 34 => tone <=b"0000000000001000";
						when 35 => tone <=b"0000000000010000";
						when 36 => tone <=b"0000000000001000";
						when 37 => tone <=b"0000000000000100";
						when 38 => tone <=b"0000000000001000";
						when 39 => tone <=b"0000000000010000";
						when 40 => tone <=b"0000000000001000";
						when 41 => tone <=b"0000000000000100";
						when 42 => tone <=b"0000000000001000";
						when 43 => tone <=b"0000000000010000";
						when 44 => tone <=b"0000000000010000";
						when 45 => tone <=b"0000000000001000";
						when 46 => tone <=b"0000000000010000";
						when 47 => tone <=b"0000010000000000";
						when 48 => tone <=b"0000001000000000";
						when 49 => tone <=b"0000000000000010";
						when 50 => tone <=b"0000000000000100";
						when 51 => tone <=b"0000000000001000";
						when 52 => tone <=b"0000000000000100";
						when 53 => tone <=b"0000000000001000";
						when 54 => tone <=b"0000001000000000";
						when 55 => tone <=b"0000000100000000";
						when 56 => tone <=b"0000000001000000";
						when 57 => tone <=b"0000000000100000";
						when 58 => tone <=b"0000000001000000";
						when 59 => tone <=b"0000000010000000";
						when others => tone <=b"0000000000000000";
					end case;
					count <= count+1;
				else
					count<=0;
				end if;
			end if;
		end if;
	end process ; -- play

	--play
	----------------------------------------------------------------------------


end architecture ; -- arch

--architecture
--------------------------------------------------------------------------------
