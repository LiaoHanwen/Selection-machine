--------------------------------------------------------------------------------
--play music
--
--input tone
--output key
--decoder
--
--integration test 10.31
--------------------------------------------------------------------------------

--------------------------------------------------------------------------------
--head

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

--head
--------------------------------------------------------------------------------

--------------------------------------------------------------------------------
--entity

entity play_music is
  port( 
  	--in
  	tone : in std_logic_vector(15 downto 0);
	
	--out
	key: out integer range 0 to 2047
  ) ;
end entity ; -- play_music

--entity
--------------------------------------------------------------------------------

--------------------------------------------------------------------------------
--architecture

architecture arch of play_music is
begin
	
	----------------------------------------------------------------------------
	--decoder

	process(tone)
		begin
			case tone is
				when "0000000000000000"  =>  key <=0;
				when "0000000000000001"  =>  key <=960;
				when "0000000000000010"  =>  key <=856;
				when "0000000000000100"  =>  key <=762;
				when "0000000000001000"  =>  key <=720;
				when "0000000000010000"  =>  key <=643;
				when "0000000000100000"  =>  key <=572;
				when "0000000001000000"  =>  key <=508;
				when "0000000010000000"  =>  key <=480;
				when "0000000100000000"  =>  key <=240;
				when "0000001000000000"  =>  key <=214;
				when "0000010000000000"  =>  key <=190;
				when "0000100000000000"  =>  key <=180;
				when "0001000000000000"  =>  key <=160;
				when "0010000000000000"  =>  key <=143;
				when "0100000000000000"  =>  key <=127;
				when "1000000000000000"  =>  key <=430;
				when others => key <=0;
				end case;
	end process ;

	--decoder
	----------------------------------------------------------------------------
	
end architecture ; -- arch

--architecture
--------------------------------------------------------------------------------